package  sobel_config_pkg;
  parameter IMAGE_ROW_SIZE    = 8;
  parameter IMAGE_COLUMN_SIZE = 8;

  parameter THRESHOLD = 100;

  parameter string INPUT_FILE_PATH    = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/lena_hex.txt";
  parameter string OUTPUT_FILE_PATH   = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/sobel_out.txt";
endpackage