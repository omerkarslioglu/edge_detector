package  sobel_config_pkg;
  localparam IMAGE_ROW_SIZE             = 256;
  localparam IMAGE_COLUMN_SIZE          = 256;
  localparam THRESHOLD                  = 100;
  localparam string INPUT_FILE_PATH     = "C:/Users/omer/github_projects/sobel/src/picha.txt";
  localparam string OUTPUT_FILE_PATH    = "C:/Users/omer/github_projects/sobel/src/matlab/sobel_out.txt";
endpackage