package  sobel_config_pkg;
  localparam IMAGE_ROW_SIZE             = 256;
  localparam IMAGE_COLUMN_SIZE          = 256;
  localparam THRESHOLD                  = 100;
  localparam string INPUT_FILE_PATH     = "<input_file_path>;
  localparam string OUTPUT_FILE_PATH    = "<output_file_path>";
endpackage