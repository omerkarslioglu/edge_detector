package  sobel_config_pkg;
  localparam IMAGE_ROW_SIZE = 256;
  localparam IMAGE_COLUMN_SIZE = 256;
  localparam THRESHOLD = 150;
  localparam string INPUT_FILE_PATH    = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/lena_hex.txt";
  localparam string OUTPUT_FILE_PATH   = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/output_test_file.txt";
endpackage