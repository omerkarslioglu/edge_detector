package  sobel_config_pkg;
  parameter IMAGE_ROW_SIZE    = 5;
  parameter IMAGE_COLUMN_SIZE = 5;

  parameter THRESHOLD = 100;

  parameter string INPUT_FILE_PATH    = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/input_test_file.txt";
  parameter string OUTPUT_FILE_PATH   = "C:/Users/omer/Desktop/YL/BirinciDonemDersler/EE562-HDLBasedDigitalDesign/sobel/src/output_test_file.txt";
endpackage